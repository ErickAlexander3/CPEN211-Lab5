//testbench for the register file
module regfile_tb()
	//testbench does not take any inputs or outputs

	
	

endmodule
