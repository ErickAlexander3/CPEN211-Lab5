module registers()

endmodule

module decoders()
endmodule

module mux()
endmodule

module ALUX ()
