//synthesizable code for the register file
module regfile()






endmodule